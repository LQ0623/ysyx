/**
  系统寄存器堆（面积优化版）
  - 去除 MuxKey，使用 case 进行译码
  - 仅为可写 CSR 建立寄存器：MTVEC、MEPC、MCAUSE
  - MSTATUS/MVENDORID/MARCHID 直接组合逻辑返回常量
  - 写入与中断处理放在同一 always 块中（irq 优先）
*/
`timescale 1ns/1ps

`define MSTATUS   12'h300
`define MTVEC     12'h305
`define MCAUSE    12'h342
`define MEPC      12'h341
`define MVENDORID 12'hF11   // 厂商 ID（Vendor ID）
`define MARCHID   12'hF12   // 架构 ID（Architecture ID）

module ysyx_24100006_CSR #(
  parameter ADDR_WIDTH = 12,
  parameter DATA_WIDTH = 32
)(
  input                       clk,
  input                       irq,
  input       [3:0]           irq_no,          // 中断号（低 8 位）
  input       [DATA_WIDTH-1:0] wdata,
  input       [ADDR_WIDTH-1:0] waddr,
  input                       wen,
  input       [ADDR_WIDTH-1:0] raddr,          // csr 指令的 31-20 位
  output reg  [DATA_WIDTH-1:0] rdata,
  output reg  [DATA_WIDTH-1:0] mtvec,
  output reg  [DATA_WIDTH-1:0] mepc
);

  // ===== 只读/常量 CSR（组合逻辑返回，不占用触发器） =====
  // 与原实现保持一致
  localparam [DATA_WIDTH-1:0] MSTATUS_CONST   = 32'h00001800; // 原代码固定写为 0x1800
  localparam [DATA_WIDTH-1:0] MVENDORID_CONST = 32'h79737978; // 'ysyx'
  localparam [DATA_WIDTH-1:0] MARCHID_CONST   = 32'd24100006; // 工程 ID

  // ===== 可写 CSR（最小集合）：MTVEC、MEPC、MCAUSE =====
  reg [3:0] mcause;

  // ===== 写入与中断处理（合并为一个时序块；irq 优先） =====
  always @(posedge clk) begin
    if (irq) begin
      // 中断到来：记录中断原因与返回地址
      mcause <= irq_no; // 高位清零，低 8 位为 irq_no
      mepc   <= wdata;                             // 与原实现一致：irq 时 mepc <- wdata
    end
    else if (wen) begin
      // 普通 CSR 写：仅允许写 MTVEC/MEPC/MCAUSE
      case (waddr)
        `MTVEC:  mtvec  <= wdata;
        `MEPC:   mepc   <= wdata;
        `MCAUSE: mcause <= wdata[3:0];
        default: ; // 其他 CSR 忽略写（MSTATUS/MVENDORID/MARCHID 为只读/常量）
      endcase
    end
  end

  // ===== CSR 读：组合译码 =====
  always @* begin
    case (raddr)
      `MSTATUS:   rdata = MSTATUS_CONST;    // 只读常量
      `MTVEC:     rdata = mtvec;            // 可写寄存器
      `MCAUSE:    rdata = { 28'b0, mcause};           // 可写寄存器
      `MEPC:      rdata = mepc;             // 可写寄存器
      `MVENDORID: rdata = MVENDORID_CONST;  // 只读常量
      `MARCHID:   rdata = MARCHID_CONST;    // 只读常量
      default:    rdata = {DATA_WIDTH{1'b0}};
    endcase
  end

`ifdef VERILATOR_SIM
import "DPI-C" function void get_csr(
	input int mstatus, 
	input int mtvec, 
	input int mcause, 
	input int mepc
);
  always @(*) begin
    get_csr(32'h00001800, mtvec, {28'b0,mcause}, mepc);
  end

`endif




endmodule
